`ifndef __DUT_REG_PKG__
`define __DUT_REG_PKG__

package dut_reg_pkg;

    `include "dut_reg_common.svh"

    `include "dut_reg_1_reg.sv"
    `include "dut_reg_2_reg.sv"
    `include "dut_reg_block.sv"

endpackage

`endif
