package uvm_hello_world_pkg;
	import uvm_pkg::*;

	`include "uvm_hello_world_test.sv"
endpackage : uvm_hello_world_pkg