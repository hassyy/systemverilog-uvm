`ifndef __SEQUENCE_COMMON__
`define __SEQUENCE_COMMON__

import uvm_pkg::*;
`include "uvm_macros.svh"

//`include "sequence_define.svh"

import image_pipe_pkg::*;
import reg_cpu_pkg::*;
import reset_pkg::*;
import dut_reg_pkg::*;

`endif
