`ifndef __RESET_DEFINE__
`define __RESET_DEFINE__

    `define RESET_RESET_ACTIVE 1'b0
    `define RESET_RESET_INACTIVE !`RESET_RESET_ACTIVE

`endif