`ifndef __TEST_PKG__
`define __TEST_PKG__

package test_pkg;

    `include "test_common.svh"

    import sequence_pkg::*;

    `include "test_lib.sv"
    `include "image_pipe_primary_test.sv"

endpackage

`endif
