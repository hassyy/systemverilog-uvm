`ifndef __DEFINE__
    `define __DEFINE__

    `define RESET_ACTIVE 0
    `define RESET_CYCLE 2
    `define CLK_PERIOD 10


`endif