`ifndef __TEST_COMMON__
`define __TEST_COMMON__

import uvm_pkg::*;
`include "uvm_macros.svh"

import image_pipe_pkg::*;
import dut_env_pkg::*;
import dut_reg_pkg::*;

// `include "test_define.svh"

`endif
