`ifndef __DUT_REG_COMMON__
`define __DUT_REG_COMMON__

import uvm_pkg::*;
`include "uvm_macros.svh"

// `include "dut_reg_define.svh"

`endif