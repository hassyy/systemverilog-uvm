`ifndef __IMAGE_PIPE_COMMON__
`define __IMAGE_PIPE_COMMON__

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "image_pipe_define.svh"

`endif
