`ifndef __TEST_COMMON__
`define __TEST_COMMON__

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "test_define.svh"

`endif
