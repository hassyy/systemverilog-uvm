`ifndef __DUT_ENV_COMMON__
`define __DUT_ENV_COMMON__

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "dut_env_define.svh"

`endif
