`ifndef __REG_CPU_COMMON__
`define __REG_CPU_COMMON__

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "reset_define.svh"

`endif