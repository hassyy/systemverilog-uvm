`ifndef __REG_CPU_REG_PREDICTOR__
`define __REG_CPU_REG_PREDICTOR__

`include "reg_cpu_common.svh"
`include "reg_cpu_data.sv"

typedef uvm_reg_predictor#(reg_cpu_data#()) reg_cpu_reg_predictor;

`endif
