`ifndef __DEFINE__
    `define __DEFINE__

    `define RESET_ACTIVE 0
    `define RESET_CYCLE 2
    `define CLK_PERIOD 10

    `define IMAGE_PIPE_DW_IN1  32
    `define IMAGE_PIPE_DW_OUT1 32


`endif