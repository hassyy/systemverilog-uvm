
`ifndef __COMMON_HEADER__
`define __COMMON_HEADER__

    import uvm_pkg::*;
    `include "uvm_macros.svh"

`endif

