`ifndef __REG_CPU_DRIVER__
    `define __REG_CPU_DRIVER__

`include "common_header.svh"
`include "define.svh"
`include "reg_cpu_data.sv"

`endif