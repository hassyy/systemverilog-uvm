`ifndef __RESET_PKG__
`define __RESET_PKG__

package reset_pkg;

    `include "reset_common.svh"

    `include "reset_transaction.sv"
    `include "reset_driver.sv"
    `include "reset_sequencer.sv"
    `include "reset_sequence.sv"

endpackage

`endif
